library verilog;
use verilog.vl_types.all;
entity Bit_sync_tb is
end Bit_sync_tb;
