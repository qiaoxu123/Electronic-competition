library verilog;
use verilog.vl_types.all;
entity tb_2011 is
end tb_2011;
