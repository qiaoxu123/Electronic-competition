module	cycle(
		//system	interface
		input			clk,
		input			rst_n,
		//sig_in	interface
		input			sig_in,
		input			sig_in1
);

//���ؼ��
reg				pulse_sig;
reg				pulse_sig1;

	



endmodule