module		

pinlv(
		//system	interface
		input					clk,
		input					rst_n,
		//sig		interface
		input					sig_in
		//user		interface
		output	reg	[31:0]		pinlv

);



endmodule