library verilog;
use verilog.vl_types.all;
entity tb_2003 is
end tb_2003;
