library verilog;
use verilog.vl_types.all;
entity hmc830_vlg_tst is
end hmc830_vlg_tst;
