library verilog;
use verilog.vl_types.all;
entity tb_uart is
end tb_uart;
