library verilog;
use verilog.vl_types.all;
entity M_sequence_tb is
end M_sequence_tb;
