library verilog;
use verilog.vl_types.all;
entity HMC830_vlg_tst is
end HMC830_vlg_tst;
