library verilog;
use verilog.vl_types.all;
entity vga_test_tb is
end vga_test_tb;
