// cpu.v

// Generated using ACDS version 13.1 162 at 2017.06.28.11:18:38

`timescale 1 ps / 1 ps
module cpu (
		input  wire        clk_clk,              //           clk.clk
		input  wire        reset_reset_n,        //         reset.reset_n
		output wire [12:0] sdram_addr,           //         sdram.addr
		output wire [1:0]  sdram_ba,             //              .ba
		output wire        sdram_cas_n,          //              .cas_n
		output wire        sdram_cke,            //              .cke
		output wire        sdram_cs_n,           //              .cs_n
		inout  wire [15:0] sdram_dq,             //              .dq
		output wire [1:0]  sdram_dqm,            //              .dqm
		output wire        sdram_ras_n,          //              .ras_n
		output wire        sdram_we_n,           //              .we_n
		input  wire        uart_rxd,             //          uart.rxd
		output wire        uart_txd,             //              .txd
		input  wire [31:0] freq_a_export,        //        freq_a.export
		input  wire [31:0] freq_b_export,        //        freq_b.export
		input  wire [31:0] freq_standard_export, // freq_standard.export
		input  wire [31:0] time_interval_export, // time_interval.export
		input  wire [31:0] duty_cycle_a_export,  //  duty_cycle_a.export
		input  wire [31:0] duty_cycle_b_export,  //  duty_cycle_b.export
		input  wire [31:0] whole_time_a_export,  //  whole_time_a.export
		input  wire [31:0] whole_time_b_export   //  whole_time_b.export
	);

	wire  [15:0] mm_interconnect_0_timer_10ms_s1_writedata;                   // mm_interconnect_0:timer_10ms_s1_writedata -> timer_10ms:writedata
	wire   [2:0] mm_interconnect_0_timer_10ms_s1_address;                     // mm_interconnect_0:timer_10ms_s1_address -> timer_10ms:address
	wire         mm_interconnect_0_timer_10ms_s1_chipselect;                  // mm_interconnect_0:timer_10ms_s1_chipselect -> timer_10ms:chipselect
	wire         mm_interconnect_0_timer_10ms_s1_write;                       // mm_interconnect_0:timer_10ms_s1_write -> timer_10ms:write_n
	wire  [15:0] mm_interconnect_0_timer_10ms_s1_readdata;                    // timer_10ms:readdata -> mm_interconnect_0:timer_10ms_s1_readdata
	wire         cpu_instruction_master_waitrequest;                          // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [27:0] cpu_instruction_master_address;                              // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                 // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire  [31:0] cpu_instruction_master_readdata;                             // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_readdatavalid;                        // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire   [1:0] mm_interconnect_0_duty_cycle_a_s1_address;                   // mm_interconnect_0:Duty_cycle_a_s1_address -> Duty_cycle_a:address
	wire  [31:0] mm_interconnect_0_duty_cycle_a_s1_readdata;                  // Duty_cycle_a:readdata -> mm_interconnect_0:Duty_cycle_a_s1_readdata
	wire   [0:0] mm_interconnect_0_sysid0_control_slave_address;              // mm_interconnect_0:sysid0_control_slave_address -> sysid0:address
	wire  [31:0] mm_interconnect_0_sysid0_control_slave_readdata;             // sysid0:readdata -> mm_interconnect_0:sysid0_control_slave_readdata
	wire   [1:0] mm_interconnect_0_freq_standard_s1_address;                  // mm_interconnect_0:Freq_standard_s1_address -> Freq_standard:address
	wire  [31:0] mm_interconnect_0_freq_standard_s1_readdata;                 // Freq_standard:readdata -> mm_interconnect_0:Freq_standard_s1_readdata
	wire  [15:0] mm_interconnect_0_uart_s1_writedata;                         // mm_interconnect_0:uart_s1_writedata -> uart:writedata
	wire   [2:0] mm_interconnect_0_uart_s1_address;                           // mm_interconnect_0:uart_s1_address -> uart:address
	wire         mm_interconnect_0_uart_s1_chipselect;                        // mm_interconnect_0:uart_s1_chipselect -> uart:chipselect
	wire         mm_interconnect_0_uart_s1_write;                             // mm_interconnect_0:uart_s1_write -> uart:write_n
	wire         mm_interconnect_0_uart_s1_read;                              // mm_interconnect_0:uart_s1_read -> uart:read_n
	wire  [15:0] mm_interconnect_0_uart_s1_readdata;                          // uart:readdata -> mm_interconnect_0:uart_s1_readdata
	wire         mm_interconnect_0_uart_s1_begintransfer;                     // mm_interconnect_0:uart_s1_begintransfer -> uart:begintransfer
	wire   [1:0] mm_interconnect_0_whole_time_b_s1_address;                   // mm_interconnect_0:Whole_time_b_s1_address -> Whole_time_b:address
	wire  [31:0] mm_interconnect_0_whole_time_b_s1_readdata;                  // Whole_time_b:readdata -> mm_interconnect_0:Whole_time_b_s1_readdata
	wire   [1:0] mm_interconnect_0_freq_a_s1_address;                         // mm_interconnect_0:Freq_a_s1_address -> Freq_a:address
	wire  [31:0] mm_interconnect_0_freq_a_s1_readdata;                        // Freq_a:readdata -> mm_interconnect_0:Freq_a_s1_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;         // cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;           // mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;             // mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;               // mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;                // mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;            // cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;         // mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;          // mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	wire         cpu_data_master_waitrequest;                                 // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire  [31:0] cpu_data_master_writedata;                                   // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [27:0] cpu_data_master_address;                                     // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire         cpu_data_master_write;                                       // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire         cpu_data_master_read;                                        // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire  [31:0] cpu_data_master_readdata;                                    // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_debugaccess;                                 // cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire         cpu_data_master_readdatavalid;                               // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire   [3:0] cpu_data_master_byteenable;                                  // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire   [1:0] mm_interconnect_0_freq_b_s1_address;                         // mm_interconnect_0:Freq_b_s1_address -> Freq_b:address
	wire  [31:0] mm_interconnect_0_freq_b_s1_readdata;                        // Freq_b:readdata -> mm_interconnect_0:Freq_b_s1_readdata
	wire   [1:0] mm_interconnect_0_whole_time_a_s1_address;                   // mm_interconnect_0:Whole_time_a_s1_address -> Whole_time_a:address
	wire  [31:0] mm_interconnect_0_whole_time_a_s1_readdata;                  // Whole_time_a:readdata -> mm_interconnect_0:Whole_time_a_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                      // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                        // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                          // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_chipselect;                       // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire         mm_interconnect_0_sdram_s1_write;                            // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire         mm_interconnect_0_sdram_s1_read;                             // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                         // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                    // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                       // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire   [1:0] mm_interconnect_0_duty_cycle_b_s1_address;                   // mm_interconnect_0:Duty_cycle_b_s1_address -> Duty_cycle_b:address
	wire  [31:0] mm_interconnect_0_duty_cycle_b_s1_readdata;                  // Duty_cycle_b:readdata -> mm_interconnect_0:Duty_cycle_b_s1_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire   [1:0] mm_interconnect_0_time_interval_s1_address;                  // mm_interconnect_0:Time_interval_s1_address -> Time_interval:address
	wire  [31:0] mm_interconnect_0_time_interval_s1_readdata;                 // Time_interval:readdata -> mm_interconnect_0:Time_interval_s1_readdata
	wire         irq_mapper_receiver0_irq;                                    // timer_10ms:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                    // uart:irq -> irq_mapper:receiver2_irq
	wire  [31:0] cpu_d_irq_irq;                                               // irq_mapper:sender_irq -> cpu:d_irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [Duty_cycle_a:reset_n, Duty_cycle_b:reset_n, Freq_a:reset_n, Freq_b:reset_n, Freq_standard:reset_n, Time_interval:reset_n, Whole_time_a:reset_n, Whole_time_b:reset_n, cpu:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset, rst_translator:in_reset, sdram:reset_n, sysid0:reset_n, timer_10ms:reset_n, uart:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]

	cpu_cpu cpu (
		.clk                                   (clk_clk),                                             //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                     //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (cpu_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (),                                                    //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	cpu_timer_10ms timer_10ms (
		.clk        (clk_clk),                                    //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            // reset.reset_n
		.address    (mm_interconnect_0_timer_10ms_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_10ms_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_10ms_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_10ms_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_10ms_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                    //   irq.irq
	);

	cpu_sdram sdram (
		.clk            (clk_clk),                                  //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	cpu_sysid0 sysid0 (
		.clock    (clk_clk),                                         //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_0_sysid0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid0_control_slave_address)   //              .address
	);

	cpu_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                     //               irq.irq
	);

	cpu_uart uart (
		.clk           (clk_clk),                                 //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address       (mm_interconnect_0_uart_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_s1_readdata),      //                    .readdata
		.dataavailable (),                                        //                    .dataavailable
		.readyfordata  (),                                        //                    .readyfordata
		.rxd           (uart_rxd),                                // external_connection.export
		.txd           (uart_txd),                                //                    .export
		.irq           (irq_mapper_receiver2_irq)                 //                 irq.irq
	);

	cpu_Freq_a freq_a (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_freq_a_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_freq_a_s1_readdata), //                    .readdata
		.in_port  (freq_a_export)                         // external_connection.export
	);

	cpu_Freq_a freq_b (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_freq_b_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_freq_b_s1_readdata), //                    .readdata
		.in_port  (freq_b_export)                         // external_connection.export
	);

	cpu_Freq_a freq_standard (
		.clk      (clk_clk),                                     //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address  (mm_interconnect_0_freq_standard_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_freq_standard_s1_readdata), //                    .readdata
		.in_port  (freq_standard_export)                         // external_connection.export
	);

	cpu_Freq_a time_interval (
		.clk      (clk_clk),                                     //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address  (mm_interconnect_0_time_interval_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_time_interval_s1_readdata), //                    .readdata
		.in_port  (time_interval_export)                         // external_connection.export
	);

	cpu_Freq_a duty_cycle_a (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_duty_cycle_a_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_duty_cycle_a_s1_readdata), //                    .readdata
		.in_port  (duty_cycle_a_export)                         // external_connection.export
	);

	cpu_Freq_a duty_cycle_b (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_duty_cycle_b_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_duty_cycle_b_s1_readdata), //                    .readdata
		.in_port  (duty_cycle_b_export)                         // external_connection.export
	);

	cpu_Freq_a whole_time_a (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_whole_time_a_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_whole_time_a_s1_readdata), //                    .readdata
		.in_port  (whole_time_a_export)                         // external_connection.export
	);

	cpu_Freq_a whole_time_b (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_whole_time_b_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_whole_time_b_s1_readdata), //                    .readdata
		.in_port  (whole_time_b_export)                         // external_connection.export
	);

	cpu_mm_interconnect_0 mm_interconnect_0 (
		.clk_100_clk_clk                           (clk_clk),                                                     //                       clk_100_clk.clk
		.cpu_reset_n_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                              // cpu_reset_n_reset_bridge_in_reset.reset
		.cpu_data_master_address                   (cpu_data_master_address),                                     //                   cpu_data_master.address
		.cpu_data_master_waitrequest               (cpu_data_master_waitrequest),                                 //                                  .waitrequest
		.cpu_data_master_byteenable                (cpu_data_master_byteenable),                                  //                                  .byteenable
		.cpu_data_master_read                      (cpu_data_master_read),                                        //                                  .read
		.cpu_data_master_readdata                  (cpu_data_master_readdata),                                    //                                  .readdata
		.cpu_data_master_readdatavalid             (cpu_data_master_readdatavalid),                               //                                  .readdatavalid
		.cpu_data_master_write                     (cpu_data_master_write),                                       //                                  .write
		.cpu_data_master_writedata                 (cpu_data_master_writedata),                                   //                                  .writedata
		.cpu_data_master_debugaccess               (cpu_data_master_debugaccess),                                 //                                  .debugaccess
		.cpu_instruction_master_address            (cpu_instruction_master_address),                              //            cpu_instruction_master.address
		.cpu_instruction_master_waitrequest        (cpu_instruction_master_waitrequest),                          //                                  .waitrequest
		.cpu_instruction_master_read               (cpu_instruction_master_read),                                 //                                  .read
		.cpu_instruction_master_readdata           (cpu_instruction_master_readdata),                             //                                  .readdata
		.cpu_instruction_master_readdatavalid      (cpu_instruction_master_readdatavalid),                        //                                  .readdatavalid
		.cpu_jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),             //             cpu_jtag_debug_module.address
		.cpu_jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),               //                                  .write
		.cpu_jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),                //                                  .read
		.cpu_jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),            //                                  .readdata
		.cpu_jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),           //                                  .writedata
		.cpu_jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),          //                                  .byteenable
		.cpu_jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),         //                                  .waitrequest
		.cpu_jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),         //                                  .debugaccess
		.Duty_cycle_a_s1_address                   (mm_interconnect_0_duty_cycle_a_s1_address),                   //                   Duty_cycle_a_s1.address
		.Duty_cycle_a_s1_readdata                  (mm_interconnect_0_duty_cycle_a_s1_readdata),                  //                                  .readdata
		.Duty_cycle_b_s1_address                   (mm_interconnect_0_duty_cycle_b_s1_address),                   //                   Duty_cycle_b_s1.address
		.Duty_cycle_b_s1_readdata                  (mm_interconnect_0_duty_cycle_b_s1_readdata),                  //                                  .readdata
		.Freq_a_s1_address                         (mm_interconnect_0_freq_a_s1_address),                         //                         Freq_a_s1.address
		.Freq_a_s1_readdata                        (mm_interconnect_0_freq_a_s1_readdata),                        //                                  .readdata
		.Freq_b_s1_address                         (mm_interconnect_0_freq_b_s1_address),                         //                         Freq_b_s1.address
		.Freq_b_s1_readdata                        (mm_interconnect_0_freq_b_s1_readdata),                        //                                  .readdata
		.Freq_standard_s1_address                  (mm_interconnect_0_freq_standard_s1_address),                  //                  Freq_standard_s1.address
		.Freq_standard_s1_readdata                 (mm_interconnect_0_freq_standard_s1_readdata),                 //                                  .readdata
		.jtag_uart_0_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //     jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                  .write
		.jtag_uart_0_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                  .read
		.jtag_uart_0_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                  .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                  .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                  .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                  .chipselect
		.sdram_s1_address                          (mm_interconnect_0_sdram_s1_address),                          //                          sdram_s1.address
		.sdram_s1_write                            (mm_interconnect_0_sdram_s1_write),                            //                                  .write
		.sdram_s1_read                             (mm_interconnect_0_sdram_s1_read),                             //                                  .read
		.sdram_s1_readdata                         (mm_interconnect_0_sdram_s1_readdata),                         //                                  .readdata
		.sdram_s1_writedata                        (mm_interconnect_0_sdram_s1_writedata),                        //                                  .writedata
		.sdram_s1_byteenable                       (mm_interconnect_0_sdram_s1_byteenable),                       //                                  .byteenable
		.sdram_s1_readdatavalid                    (mm_interconnect_0_sdram_s1_readdatavalid),                    //                                  .readdatavalid
		.sdram_s1_waitrequest                      (mm_interconnect_0_sdram_s1_waitrequest),                      //                                  .waitrequest
		.sdram_s1_chipselect                       (mm_interconnect_0_sdram_s1_chipselect),                       //                                  .chipselect
		.sysid0_control_slave_address              (mm_interconnect_0_sysid0_control_slave_address),              //              sysid0_control_slave.address
		.sysid0_control_slave_readdata             (mm_interconnect_0_sysid0_control_slave_readdata),             //                                  .readdata
		.Time_interval_s1_address                  (mm_interconnect_0_time_interval_s1_address),                  //                  Time_interval_s1.address
		.Time_interval_s1_readdata                 (mm_interconnect_0_time_interval_s1_readdata),                 //                                  .readdata
		.timer_10ms_s1_address                     (mm_interconnect_0_timer_10ms_s1_address),                     //                     timer_10ms_s1.address
		.timer_10ms_s1_write                       (mm_interconnect_0_timer_10ms_s1_write),                       //                                  .write
		.timer_10ms_s1_readdata                    (mm_interconnect_0_timer_10ms_s1_readdata),                    //                                  .readdata
		.timer_10ms_s1_writedata                   (mm_interconnect_0_timer_10ms_s1_writedata),                   //                                  .writedata
		.timer_10ms_s1_chipselect                  (mm_interconnect_0_timer_10ms_s1_chipselect),                  //                                  .chipselect
		.uart_s1_address                           (mm_interconnect_0_uart_s1_address),                           //                           uart_s1.address
		.uart_s1_write                             (mm_interconnect_0_uart_s1_write),                             //                                  .write
		.uart_s1_read                              (mm_interconnect_0_uart_s1_read),                              //                                  .read
		.uart_s1_readdata                          (mm_interconnect_0_uart_s1_readdata),                          //                                  .readdata
		.uart_s1_writedata                         (mm_interconnect_0_uart_s1_writedata),                         //                                  .writedata
		.uart_s1_begintransfer                     (mm_interconnect_0_uart_s1_begintransfer),                     //                                  .begintransfer
		.uart_s1_chipselect                        (mm_interconnect_0_uart_s1_chipselect),                        //                                  .chipselect
		.Whole_time_a_s1_address                   (mm_interconnect_0_whole_time_a_s1_address),                   //                   Whole_time_a_s1.address
		.Whole_time_a_s1_readdata                  (mm_interconnect_0_whole_time_a_s1_readdata),                  //                                  .readdata
		.Whole_time_b_s1_address                   (mm_interconnect_0_whole_time_b_s1_address),                   //                   Whole_time_b_s1.address
		.Whole_time_b_s1_readdata                  (mm_interconnect_0_whole_time_b_s1_readdata)                   //                                  .readdata
	);

	cpu_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (cpu_d_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
