library verilog;
use verilog.vl_types.all;
entity Digital_Freq_top_tb is
end Digital_Freq_top_tb;
