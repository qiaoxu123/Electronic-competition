library verilog;
use verilog.vl_types.all;
entity tb_2007 is
end tb_2007;
